library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package duty_cycle_pkg is
        type duty_array is array(natural range <>) of std_logic_vector;
end package;


package body duty_cycle_pkg is 

end duty_cycle_pkg; 